** sch_path: /home/thanhtung/projects/inverter/xschem/New folder/dls_nand.sch
**.subckt dls_nand
XM1 Vout Vin1 net1 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
V1 VDD GND 0.8
.save i(v1)
Vin Vin1 GND pulse( 0 0.8 0 0 0 5 10)
.save i(vin)
XM5 net1 Vin2 net2 GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 Vout Vin1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vout Vin2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 VDD Vout VDD GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 GND Vout net2 GND sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
Vin1 Vin2 GND pulse( 0.8 0 2.5 0 0 5 10)
.save i(vin1)
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/thanhtung/eda/unic-cass/share/pdk/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/thanhtung/eda/unic-cass/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/thanhtung/eda/unic-cass/share/pdk/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/thanhtung/eda/unic-cass/share/pdk/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice



.save all
.control
tran 0.1 50
meas tran curr_avg avg v1#branch from=0s to=50s
let P=curr_avg*0.8
print P>>Power_dls.txt
set color0=white
set colot1=black
set color2=purple
set xbrushwidth=5
plot Vin1+2 Vin2+1 Vout+0
.endc



**** end user architecture code
**.ends
.GLOBAL GND
.GLOBAL VDD
.end
